module tile_tb();




endmodule